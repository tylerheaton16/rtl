module PulseSynchronizer (
  input clkA, clkB,
  input resetn,
  input sig1,
  output wire sig_sync
);

endmodule
